// Lucas Lemos - llemos@hmc.edu - 9/2/2025
// Tests the top level module of the lab2_ll_two_displays project.
// Tests that the LED count adder computes the right value based on the two input switches
// and the switch select mux properly oscillates according to the divided clock.

// Questa requires a timescale 
`timescale 1 ms / 1 ms

module lab_2_ll_tb;
	// DUT logic
	logic [3:0] switch1, switch2; // input
	logic       reset_p34;        // input
	logic       clk_div_p2;       // output
	logic [4:0] led_cnt;          // output
	logic [6:0] seg;              // output
	
	// Testing logic unique to this DUT	
	logic [6:0] seg_expected1, seg_expected2;
	logic [4:0] led_expected;
	
	// General testbench logic	
	//logic        clk;
	logic [31:0] vectornum;            // index value of test vectors 
	logic [31:0] errors;               // number of errors
	logic [31:0] testvectors[10000:0]; // create space for 10,000 32-bit wide test vectors
	
	// Instantiate device under test	
	lab2_ll_two_displays DUT(
		.switch1    ( switch1 ),    // input [3:0]
		.switch2    ( switch2 ),    // input [3:0]
		.reset_p34  ( reset_p34 ),  // input
		.clk_div_p2 ( clk_div_p2 ), // output
		.led_cnt    ( led_cnt ),    // output [4:0]
		.seg        ( seg )        // output [6:0]
	);
		/*
	// Generate test clock	
	always
		begin
			clk=1; #5; clk=0; #5;
		end 
	*/
	// Begin test by loading vectors & pulsing reset
		initial
		begin
			$readmemb("lab2_ll_vectors.tv", testvectors);
			vectornum = 0; errors = 0; reset_p34 = 0; #12; reset_p34 = 1;
		end
	
	// Load next test vector
	always @(posedge clk_div_p2) // was clk
		begin
			#1; {switch1, switch2, seg_expected1, seg_expected2, led_expected} = testvectors[vectornum];
		end //^ THAT MIGHT NEED TO BE #2 FOR TEST VECTORS TO LOAD PROPERLY
	
	
	// Check seg outputs and led_cnt output against switch 1 & 2 inputs
	always @(posedge clk_div_p2) begin
		if (reset_p34) begin  // remember-- reset is active low
			/* // The automatic error correction is still buggy, but I can visually verify that the sim is working -- except the weird transition points on seg makes me think it is still broken (maybe has to do with how vector loading is delayed by #1?)
			// Check both seg outputs
			if (seg == seg_expected1) begin
				#1; assert(seg == seg_expected2) else begin // THAT #1 MIGHT NEED TO BE WAY BIGGER
					$error("Error: one of two segs failed.");
					$display("switch1: %b, switch2: %b, seg: %b, seg_expected1: %b, seg_expected2: %b", switch1, switch2, seg, seg_expected1, seg_expected2);
					errors = errors + 1;
				end
			end
			else if (seg == seg_expected2) begin
				#1; assert(seg == seg_expected1) else begin // THAT #1 MIGHT NEED TO BE WAY BIGGER
					$error("Error: one of two segs failed.");
					$display("switch1: %b, switch2: %b, seg: %b, seg_expected1: %b, seg_expected2: %b", switch1, switch2, seg, seg_expected1, seg_expected2);
					errors = errors + 1;
				end
			end
			else begin
				$error("Both segs failed.");
				$display("switch1: %b, switch2: %b, seg: %b, seg_expected1: %b, seg_expected2: %b", switch1, switch2, seg, seg_expected1, seg_expected2);
				errors = errors + 1;
			end
			
			// Check led_cnt
			assert(led_cnt == led_expected) else begin
				$error("LED count failed.");
				$display("switch1: %b, switch2: %b, led_cnt: %b, led_expected: %b", switch1, switch2, led_cnt, led_expected);
			end
			*/
		vectornum = vectornum + 1;
		
		// Check if simulation has ended
		if (testvectors[vectornum] === 32'bx) begin
				$display("%d tests completed with %d errors", vectornum, errors);
				$stop;	// End the simulation
			end
		end
	end
endmodule

	/*
	// check results on falling edge of clk
always @(negedge clk)
 if (~reset) begin // skip during reset
 if ({la, lb, lc, ra, rb, rc} !== expected) begin // check result
 $display("Error: inputs = %b", {left, right});
 $display(" outputs = %b %b %b %b %b %b (%b expected)",
 la, lb, lc, ra, rb, rc, expected);
 errors = errors + 1;
 end
 vectornum = vectornum + 1;
 if (testvectors[vectornum] === 8'bx) begin
 $display("%d tests completed with %d errors", vectornum, errors);
 $stop;
 end
 end
endmodule 
*/
	
