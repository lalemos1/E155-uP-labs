// Lucas Lemos - llemos@hmc.edu - 9/15/2025
// This top level module



// DON'T USE SYNCHRONIZER FOR NOW--GET MVP WORKING